module ggui
import gx

pub struct CatppuchinMocha {
pub:
	crust	   gx.Color = gx.Color{17, 17, 27, 255}
	mantle	   gx.Color = gx.Color{24, 24, 37, 255}
	base	   gx.Color = gx.Color{30, 30, 46, 255}
	surface0   gx.Color = gx.Color{49, 50, 68, 255}
	surface1   gx.Color = gx.Color{69, 71, 90, 255}
	surface2   gx.Color = gx.Color{88, 91, 112, 255}
	overlay0   gx.Color = gx.Color{108, 112, 134, 255}
	overlay1   gx.Color = gx.Color{127, 132, 156, 255}
	overlay2   gx.Color = gx.Color{147, 153, 178, 255}
	subtext0   gx.Color = gx.Color{166, 173, 200, 255}
	subtext1   gx.Color = gx.Color{186, 194, 222, 255}
	text	   gx.Color = gx.Color{205, 214, 244, 255}
	lavender   gx.Color = gx.Color{180, 190, 254, 255}
	blue	   gx.Color = gx.Color{137, 180, 250, 255}
	sapphire   gx.Color = gx.Color{116, 199, 236, 255}
	sky		   gx.Color = gx.Color{137, 220, 235, 255}
	teal	   gx.Color = gx.Color{148, 227, 213, 255}
	green	   gx.Color = gx.Color{166, 214, 161, 255}
	yellow	   gx.Color = gx.Color{249, 226, 175, 255}
	peach	   gx.Color = gx.Color{250, 179, 135, 255}
	maroon	   gx.Color = gx.Color{235, 160, 172, 255}
	red		   gx.Color = gx.Color{243, 139, 168, 255}
	mauve	   gx.Color = gx.Color{203, 166, 247, 255}
	pink	   gx.Color = gx.Color{245, 194, 231, 255}
	flamingo   gx.Color = gx.Color{242, 205, 205, 255}
	rosewater  gx.Color = gx.Color{245, 224, 220, 255}
}

pub struct CatppuchinFrappe {
pub:
	crust	   gx.Color = gx.Color{35, 38, 52, 255}
	mantle	   gx.Color = gx.Color{41, 44, 60, 255}
	base	   gx.Color = gx.Color{48, 52, 70, 255}
	surface0   gx.Color = gx.Color{65, 69, 89, 255}
	surface1   gx.Color = gx.Color{81, 87, 109, 255}
	surface2   gx.Color = gx.Color{98, 104, 128, 255}
	overlay0   gx.Color = gx.Color{115, 121, 148, 255}
	overlay1   gx.Color = gx.Color{131, 139, 167, 255}
	overlay2   gx.Color = gx.Color{148, 156, 187, 255}
	subtext0   gx.Color = gx.Color{165, 173, 206, 255}
	subtext1   gx.Color = gx.Color{181, 191, 226, 255}
	text	   gx.Color = gx.Color{198, 208, 245, 255}
	lavender   gx.Color = gx.Color{186, 187, 241, 255}
	blue	   gx.Color = gx.Color{140, 170, 238, 255}
	sapphire   gx.Color = gx.Color{133, 193, 220, 255}
	sky		   gx.Color = gx.Color{153, 209, 219, 255}
	teal	   gx.Color = gx.Color{129, 200, 190, 255}
	green	   gx.Color = gx.Color{166, 209, 137, 255}
	yellow	   gx.Color = gx.Color{229, 200, 144, 255}
	peach	   gx.Color = gx.Color{239, 159, 118, 255}
	maroon	   gx.Color = gx.Color{234, 153, 156, 255}
	red		   gx.Color = gx.Color{231, 130, 132, 255}
	mauve	   gx.Color = gx.Color{202, 158, 230, 255}
	pink	   gx.Color = gx.Color{244, 184, 228, 255}
	flamingo   gx.Color = gx.Color{238, 190, 190, 255}
	rosewater  gx.Color = gx.Color{242, 213, 207, 255}
}

pub struct CatppuchinMacchiato {
pub:
	crust	   gx.Color = gx.Color{24, 25, 38, 255}
	mantle	   gx.Color = gx.Color{30, 32, 48, 255}
	base	   gx.Color = gx.Color{36, 39, 58, 255}
	surface0   gx.Color = gx.Color{54, 58, 79, 255}
	surface1   gx.Color = gx.Color{73, 77, 100, 255}
	surface2   gx.Color = gx.Color{91, 96, 120, 255}
	overlay0   gx.Color = gx.Color{110, 115, 141, 255}
	overlay1   gx.Color = gx.Color{128, 135, 162, 255}
	overlay2   gx.Color = gx.Color{147, 154, 183, 255}
	subtext0   gx.Color = gx.Color{165, 173, 203, 255}
	subtext1   gx.Color = gx.Color{184, 192, 224, 255}
	text	   gx.Color = gx.Color{202, 211, 245, 255}
	lavender   gx.Color = gx.Color{183, 189, 248, 255}
	blue	   gx.Color = gx.Color{138, 173, 244, 255}
	sapphire   gx.Color = gx.Color{125, 196, 228, 255}
	sky		   gx.Color = gx.Color{145, 215, 227, 255}
	teal	   gx.Color = gx.Color{139, 213, 202, 255}
	green	   gx.Color = gx.Color{166, 218, 149, 255}
	yellow	   gx.Color = gx.Color{238, 212, 159, 255}
	peach	   gx.Color = gx.Color{245, 169, 127, 255}
	maroon	   gx.Color = gx.Color{238, 153, 160, 255}
	red		   gx.Color = gx.Color{237, 135, 150, 255}
	mauve	   gx.Color = gx.Color{198, 160, 246, 255}
	pink	   gx.Color = gx.Color{245, 189, 230, 255}
	flamingo   gx.Color = gx.Color{240, 198, 198, 255}
	rosewater  gx.Color = gx.Color{244, 219, 214, 255}
}

pub struct CatppuchinLatte {
pub:
	crust	   gx.Color = gx.Color{220, 224, 232, 255}
	mantle	   gx.Color = gx.Color{230, 233, 239, 255}
	base	   gx.Color = gx.Color{239, 241, 245, 255}
	surface0   gx.Color = gx.Color{204, 208, 218, 255}
	surface1   gx.Color = gx.Color{188, 192, 204, 255}
	surface2   gx.Color = gx.Color{172, 176, 190, 255}
	overlay0   gx.Color = gx.Color{156, 160, 176, 255}
	overlay1   gx.Color = gx.Color{140, 143, 161, 255}
	overlay2   gx.Color = gx.Color{124, 127, 147, 255}
	subtext0   gx.Color = gx.Color{108, 111, 133, 255}
	subtext1   gx.Color = gx.Color{92, 95, 119, 255}
	text	   gx.Color = gx.Color{76, 79, 105, 255}
	lavender   gx.Color = gx.Color{114, 135, 253, 255}
	blue	   gx.Color = gx.Color{30, 102, 245, 255}
	sapphire   gx.Color = gx.Color{32, 159, 181, 255}
	sky		   gx.Color = gx.Color{4, 165, 229, 255}
	teal	   gx.Color = gx.Color{23, 146, 153, 255}
	green	   gx.Color = gx.Color{64, 160, 43, 255}
	yellow	   gx.Color = gx.Color{223, 142, 29, 255}
	peach	   gx.Color = gx.Color{254, 100, 11, 255}
	maroon	   gx.Color = gx.Color{230, 69, 83, 255}
	red		   gx.Color = gx.Color{210, 15, 57, 255}
	mauve	   gx.Color = gx.Color{136, 57, 239, 255}
	pink	   gx.Color = gx.Color{234, 118, 203, 255}
	flamingo   gx.Color = gx.Color{221, 120, 120, 255}
	rosewater  gx.Color = gx.Color{220, 138, 120, 255}
}

pub interface Clickable {
mut:
	id int
	x f32
	y f32
	shape Area
	click_func fn (mut main Gui, mut parent Gui)
	render(mut g Gui, x_offset f32, y_offset f32)
}

pub interface Area {
mut:
	width f32
	height f32
	relative_pos Pos
}

fn (a Area) offset() (f32, f32) {
	return match a.relative_pos {
		.center {-a.width/2, -a.height/2}
		.right {0, -a.height/2}
		.left {-a.width, -a.height/2}
		.top {-a.width/2, 0}
		.bottom {-a.width/2, a.height}
		.top_right {0, 0}
		.top_left {-a.width, 0}
		.bottom_right {0, a.height}
		.bottom_left {a.height, a.width}
	}
}

pub fn (a Area) render(mut g Gui, x_offset f32, y_offset f32, color gx.Color) {
	mut x_coo := x_offset
	mut y_coo := y_offset
	match a.relative_pos {
		.center {
			x_coo -= a.width/2
			y_coo -= a.height/2
		}
		.right {y_coo -= a.height/2}
		.left {
			x_coo -= a.width
			y_coo -= a.height/2
		}
		.top {x_coo -= a.width/2}
		.bottom {
			x_coo -= a.width/2
			y_coo += a.height
		}
		.top_right {}
		.top_left {
			x_coo -= a.width
		}
		.bottom_right {
			y_coo += a.height
		}
		.bottom_left {
			y_coo += a.height
			x_coo += a.width
		}
	}
	match a {
		RoundedShape {g.gg.draw_rounded_rect_filled(x_coo, y_coo, a.width, a.height, a.rounded, color)}
		else {g.gg.draw_rect_filled(x_coo, y_coo, a.width, a.height, color)}
	}
}

pub interface Element {
mut:
	id int
	x f32
	y f32
	render(mut g Gui, x_offset f32, y_offset f32)
}

pub enum Pos {
	center
	right
	left
	top
	bottom
	top_right
	top_left
	bottom_right
	bottom_left
}

pub struct RoundedShape {
pub mut:
	width f32
	height f32
	rounded int
	relative_pos Pos
}

pub struct Shape {
pub mut:
	width f32
	height f32
	relative_pos Pos
}